`timescale 1ns/1ns
module led_test_tb;
reg clk;
reg rst_n;
wire[3:0] led;
initial
begin
	clk = 1'b0;
	rst_n = 1'b0;
	#100 rst_n = 1'b1;	
end
always#10 clk = ~clk;//50Mhz
led_test dut
(
	.clk           (clk),// ������������ʱ��: 50Mhz
	.rst_n         (rst_n),// �����������븴λ����
	.led           (led)// ���LED��,���ڿ��ƿ��������ĸ�LED(LED0~LED3)
);
endmodule 